----------------------------------------------------------------------------------
-- Engineer: Donny Percivalle
--
-- Create Date:    21:15:06 01/17/2013
-- Description:    Clock divider to drive 4-digit 7-segment display.
--                 Referenced from Bryan Mealey, Associate Professor at
--                 Cal Poly SLO.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity clk_div is
   Port (  clk : in std_logic;
          sclk : out std_logic);
end clk_div;

architecture my_clk_div of clk_div is
   constant max_count : integer := (2200);
       signal tmp_clk : std_logic := '0';
   begin
   my_div: process (clk,tmp_clk)
      variable div_cnt : integer := 0;
      begin
         if (rising_edge(clk)) then
            if (div_cnt = MAX_COUNT) then
               tmp_clk <= not tmp_clk;
                div_cnt := 0;
            else
               div_cnt := div_cnt + 1;
            end if;
         end if;
      sclk <= tmp_clk;
   end process my_div;
end my_clk_div;